// Модуль, описывающий функцию F (вариант 33) на поведенческом уровне
module lab2_behavioral(
    input  X, Y, Z, K, L, N, // Входные сигналы
    output F                 // Выходной сигнал
    );
 
    // Прямое описание функции с использованием операторов Verilog
    // ~ : НЕ (NOT)
    // | : ИЛИ (OR)
    // ^ : Исключающее ИЛИ (XOR)
    assign F = ((~X | ~Y) ^ Z) ^ (~(K ^ ~L ^ ~N));
 
endmodule